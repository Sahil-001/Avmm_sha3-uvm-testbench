`include "sha3_top.sv"
`include "sha3_seq_item.sv"
`include "avl_seq_item.sv"
`include "sha3_sequencer.sv"
`include "sha3_sequence.sv"
`include "avl_sequencer.sv"
`include "interface.sv"
`include "avl_driver.sv"
`include "sha3_avl_sequence2.sv"
`include "sha3_monitor2.sv"
`include "avl_agent.sv"
`include "sha3_agent.sv"
`include "sha3_env.sv"
`include "sha3_scoreboard.sv"
`include "../../src/rtl/sha3.v"
`include "../../src/rtl/avalon_sha3_wrapper.v"
`include "../../src/rtl/sha3_wrapper.v"
`include "random_test_parameterized.sv"
`include "random_test.sv"
